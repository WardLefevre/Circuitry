versterker
Vcc	1	0	12
Vbb	2	0	AC 0.001
C1	2	3	4u
R1	1	3	14997
R2	3	0	19706
Rc	1	4	750
Rg	5	6	75
Re	6	0	750
Ce	6	0	42u
Q1	4	3	5	BC547B
C2	4	7	42u
R12	1	7	14997
R22	7	0	19706
Rc2	1	8	750
Rg2	9	10	50
Re2	10	0	750
Ce2	10	0	42u
Q12	8	7	9	BC547B
Qbu	1	8	11	BC547B
Rbu	11	0	1k
Cbu	11	12	42u
Rl	12	0	150

.MODEL BC547B NPN(IS=2.39E-14 ISE=3.545E-15 ISC=6.272E-14 XTI=3
+ BF=294 BR=7.946 IKF=0.1357 IKR=0.1144 XTB=1.5
+ VAF=63.2 VAR=25.9 VJE=0.65 VJC=0.3997
+ RE=0.4683 RC=0.85 RB=1 RBM=1 IRB=1E-06
+ CJE=1.358E-11 CJC=3.728E-12 XCJC=0.6193 FC=0.9579
+ NF=1.008 NR=1.004 NE=1.541 NC=1.243 MJE=0.3279 MJC=0.2955
+ TF=4.391E-10 TR=1E-32 PTF=0 ITF=0.7495 VTF=2.643 XTF=120
+ EG=1.11 KF=1E-9 AF=1)
*.tran 1ns 1ms
.AC DEC 1000	3	300k
.PROBE
.END