butt
V1	1	0	AC	1
R0	1	2	50
L2	2	3	15.92n
L4	3	4	29.91n
L6	4	5	29.91n
L8	5	6	15.92n
R10	6	0	50
C1	2	0	2.21p
C3	3	0	9.75p
C5	4	0	12.73p
C7	5	0	9.75p
C9	6	0	2.21p
.AC DEC 100	100MEG	1000MEG
.PROBE
.END