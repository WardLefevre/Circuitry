buttstrip
V1	1	0	AC	1
R0	1	2	50
T1	2	0	3	0	Z0=10	F=500MEG	NL=0.0110
T2	3	0	4	0	Z0=100	F=500MEG	NL=0.0796
T3	4	0	5	0	Z0=10	F=500MEG	NL=0.0487
T4	5	0	6	0	Z0=100	F=500MEG	NL=0.1495
T5	6	0	7	0	Z0=10	F=500MEG	NL=0.0636
T6	7	0	8	0	Z0=100	F=500MEG	NL=0.1495
T7	8	0	9	0	Z0=10	F=500MEG	NL=0.0487
T8	9	0	10	0	Z0=100	F=500MEG	NL=0.0796
T9	10	0	11	0	Z0=10	F=500MEG	NL=0.0101
R10	11	0	50
.AC DEC 100	10MEG	1000MEG
.PROBE
.END